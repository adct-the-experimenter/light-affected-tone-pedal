.title KiCad schematic
.include "/usr/home/computerplayer/Circuits/spice-models/lm358.lib"
VCC1 vcc 0 dc 9
RF1 IN1- OUT1 10k
RG1 IN1- 0 1k
Rpole1 vin IN1+ 10k
Cpole1 IN1+ 0 1u
Vsignal1 vin 0 dc 0 ac 1 sin(0 0.1 50)
XU1 IN1+ IN1- OUT1 vcc 0 LMX58_LM2904
.end
